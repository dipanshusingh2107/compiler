PRINT 5+10*3
PRINT "Hellooo World"
PRINT -12 * +5
PRINT "THIS LANGUAGE IS SV" 