PRINT 123 * 23 / 24 + 13 - 45
PRINT "Helllo world"