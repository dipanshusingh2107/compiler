PRINT 2323 + 32 / 3 * 4 + 43 - 23
PRINT "Helllo world"